module boundingBox(input logic clk, input logic rst_n,
            input logic en, output logic rdy,
            output logic [7:0] addr, output logic [7:0] wrdata, output logic wren,
            output logic[10:0] xMin, output logic[10:0] xMax,
            output logic[10:0] yMin, output logic[10:0] yMax);









, 


