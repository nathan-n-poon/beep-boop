module cropping
(

);